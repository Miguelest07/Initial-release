module Commando_Inicial (
	input i_clk,
	output o_Global_Enable
);
endmodule